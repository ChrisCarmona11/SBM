library IEEE ;
use IEEE.STD_LOGIC_1164.all ;

package	constants is
	type TPicoType is ( pbtI, pbtII, pbt3, pbtS ) ;
	constant PicoType : TPicoType := pbt3 ;
	function ADDRSIZE return natural ;
	function INSTSIZE return natural ;
	function JADDRSIZE return natural ;
	function JDATASIZE return natural ;
end package ;

package body constants is
	function ADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 10 ;
		when pbt3 => return 10 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function INSTSIZE return natural is 
	begin
		case PicoType is
		when pbtI => return 16 ;
		when pbtII => return 18 ;
		when pbt3 => return 18 ;
		when pbtS => return 18 ;
		end case ;
	end ;
	function JADDRSIZE return natural is
	begin
		case PicoType is
		when pbtI => return 9 ;
		when pbtII => return 11 ;
		when pbt3 => return 11 ;
		when pbtS => return 10 ;
		end case ;
	end ;
	function JDATASIZE return natural is
	begin
		case PicoType is
		when pbtI => return 8 ;
		when pbtII => return 9 ;
		when pbt3 => return 9 ;
		when pbtS => return 20 ;
		end case ;
	end ;
end package body ;


library IEEE ;
use IEEE.STD_LOGIC_1164.all ;
use IEEE.STD_LOGIC_ARITH.all ;
use IEEE.STD_LOGIC_UNSIGNED.all ;

library unisim ;
use unisim.vcomponents.all ;

use constants.all;

entity ROM_KCPSM3 is
    port ( 
        clk : in std_logic ;
        reset : out std_logic ;
        address : in std_logic_vector( ADDRSIZE - 1 downto 0 ) ;
        instruction : out std_logic_vector( INSTSIZE - 1 downto 0 )
    ) ;
end entity ROM_KCPSM3 ;

architecture mix of ROM_KCPSM3 is
    component jtag_shifter is
        port ( 
			clk : in std_logic ;
			user1 : out std_logic ;
            write : out std_logic ;
            addr : out std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
            data : out std_logic_vector( JDATASIZE - 1 downto 0 )
        ) ;
    end component ;

    signal jaddr : std_logic_vector( JADDRSIZE - 1 downto 0 ) ;
    signal jdata : std_logic_vector( JDATASIZE - 1 downto 0 ) ;
    signal juser1 : std_logic ;
    signal jwrite : std_logic ;

    attribute INIT_00 : string ;
    attribute INIT_01 : string ;
    attribute INIT_02 : string ;
    attribute INIT_03 : string ;
    attribute INIT_04 : string ;
    attribute INIT_05 : string ;
    attribute INIT_06 : string ;
    attribute INIT_07 : string ;
    attribute INIT_08 : string ;
    attribute INIT_09 : string ;
    attribute INIT_0A : string ;
    attribute INIT_0B : string ;
    attribute INIT_0C : string ;
    attribute INIT_0D : string ;
    attribute INIT_0E : string ;
    attribute INIT_0F : string ;
    attribute INIT_10 : string ;
    attribute INIT_11 : string ;
    attribute INIT_12 : string ;
    attribute INIT_13 : string ;
    attribute INIT_14 : string ;
    attribute INIT_15 : string ;
    attribute INIT_16 : string ;
    attribute INIT_17 : string ;
    attribute INIT_18 : string ;
    attribute INIT_19 : string ;
    attribute INIT_1A : string ;
    attribute INIT_1B : string ;
    attribute INIT_1C : string ;
    attribute INIT_1D : string ;
    attribute INIT_1E : string ;
    attribute INIT_1F : string ;
    attribute INIT_20 : string ;
    attribute INIT_21 : string ;
    attribute INIT_22 : string ;
    attribute INIT_23 : string ;
    attribute INIT_24 : string ;
    attribute INIT_25 : string ;
    attribute INIT_26 : string ;
    attribute INIT_27 : string ;
    attribute INIT_28 : string ;
    attribute INIT_29 : string ;
    attribute INIT_2A : string ;
    attribute INIT_2B : string ;
    attribute INIT_2C : string ;
    attribute INIT_2D : string ;
    attribute INIT_2E : string ;
    attribute INIT_2F : string ;
    attribute INIT_30 : string ;
    attribute INIT_31 : string ;
    attribute INIT_32 : string ;
    attribute INIT_33 : string ;
    attribute INIT_34 : string ;
    attribute INIT_35 : string ;
    attribute INIT_36 : string ;
    attribute INIT_37 : string ;
    attribute INIT_38 : string ;
    attribute INIT_39 : string ;
    attribute INIT_3A : string ;
    attribute INIT_3B : string ;
    attribute INIT_3C : string ;
    attribute INIT_3D : string ;
    attribute INIT_3E : string ;
    attribute INIT_3F : string ;
    attribute INITP_00 : string ;
    attribute INITP_01 : string ;
    attribute INITP_02 : string ;
    attribute INITP_03 : string ;
    attribute INITP_04 : string ;
    attribute INITP_05 : string ;
    attribute INITP_06 : string ;
    attribute INITP_07 : string ;
begin
	I18 : if (PicoType = pbtII) or (PicoType = pbt3) generate
	    attribute INIT_00 of bram : label is "BFE00F02147DBFE00F01C0010137020003000D000E00CF04CF01CF00CF070F00" ;
	    attribute INIT_01 of bram : label is "1F705066EF481F70505FEF4C1F70505FEF6C1F70AEFD400B149ABFE00F041415" ;
	    attribute INIT_02 of bram : label is "EF721F70504CEF531F70504CEF731F705047EF411F705047EF611F705066EF68" ;
	    attribute INIT_03 of bram : label is "506BEF541F70506BEF741F70505BEF441F70505BEF641F705051EF521F705051" ;
	    attribute INIT_04 of bram : label is "00B700BB13F00186A00000B700BB12F00186A000506FEF581F70506FEF781F70" ;
	    attribute INIT_05 of bram : label is "0186A00000B700FF00BBA00000B700DB00A700A3CF040F01C202C30300BBA000" ;
	    attribute INIT_06 of bram : label is "00BBA00000B7012600BBA00000B700BB11F00186A00000B700C300BBCE0410F0" ;
	    attribute INIT_07 of bram : label is "DFF01FD0AEFEA000547ACF010F05A00000B70169CF070F000079CF070F01014A" ;
	    attribute INIT_08 of bram : label is "1AC05491EF031FD0409219C0548CEF021FD0409218C05487EF01409217C05483" ;
	    attribute INIT_09 of bram : label is "0F03C101C000C202C303AEFBA00000B70D00CE02B400FFC00F0D8D010DFF4092" ;
	    attribute INIT_0A of bram : label is "54ADAF024F0414F0A000CF040F0041024001A00050A3AF014F0040A900A3CF04" ;
	    attribute INIT_0B of bram : label is "00AC0F6B00AC0F4F00B2A00000AC0F3E00B2A00000AC0F0A00AC0F0DA000C405" ;
	    attribute INIT_0C of bram : label is "00AC0F2000F31F0000F31F1000AC0F2000AC0F7200AC0F5700B2A00000AC0F21" ;
	    attribute INIT_0D of bram : label is "00AC0F6400AC0F5200B2A00000F31F2000F31F3000AC0F2000AC0F7400AC0F61" ;
	    attribute INIT_0E of bram : label is "00F31F3000AC0F2000AC0F7400AC0F6100AC0F2000F31F0000F31F1000AC0F20" ;
	    attribute INIT_0F of bram : label is "00B2A00000AC019CAF0F1F5000AC019C0F0E0F0E0F0E0F0E15F0A00000F31F20" ;
	    attribute INIT_10 of bram : label is "00F31F3000AC0F2000AC0F3D00AC0F2000AC0F7200AC0F6400AC0F6400AC0F41" ;
	    attribute INIT_11 of bram : label is "0F2000AC0F3D00AC0F2000AC0F6100AC0F7400AC0F6100AC0F4400B200F31F20" ;
	    attribute INIT_12 of bram : label is "0F7300AC0F6900AC0F2000AC1F9000AC1F8000B2A00000F31F0000F31F1000AC" ;
	    attribute INIT_13 of bram : label is "00AC0F5200AC0F4500AC0F5000AC0F4100B2A00000AC8F30018600AC0F2000AC" ;
	    attribute INIT_14 of bram : label is "00AC0F6600AC0F6F00AC0F53A00000B700AC0F3100AC0F3100AC0F2000AC0F54" ;
	    attribute INIT_15 of bram : label is "00AC0F2000AC0F7400AC0F6500AC0F7300AC0F6500AC0F5200AC0F2000AC0F74" ;
	    attribute INIT_16 of bram : label is "0F7400AC0F6600AC0F6F00AC0F53A00000AC0F6800AC0F6700AC0F6900AC0F48" ;
	    attribute INIT_17 of bram : label is "0F4C00AC0F2000AC0F7400AC0F6500AC0F7300AC0F6500AC0F5200AC0F2000AC" ;
	    attribute INIT_18 of bram : label is "5193B880A80FA90F19F001951F9018F001951F80A00000AC0F7700AC0F6F00AC" ;
	    attribute INIT_19 of bram : label is "8F305DA1C40A14F0A000CF37A000CF305D9AC44014F0A0001F90418EC8018910" ;
	    attribute INIT_1A of bram : label is "1FC04C0316F0A00000B700BB55A4850100AC8F301F5000B205EAA0008F37A000" ;
	    attribute INIT_1B of bram : label is "00000000000000000000000000000000000000000000000080011F600E0100AC" ;
	    attribute INIT_1C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_1F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_20 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_21 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_22 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_23 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_24 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_25 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_26 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_27 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_28 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_29 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_2F of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_30 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_31 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_32 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_33 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_34 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_35 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_36 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_37 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_38 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_39 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3A of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3B of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3C of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3D of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3E of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INIT_3F of bram : label is "41AD000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_00 of bram : label is "02D2F8E3EFEF3BF0EFEFF8AEF3BCEC30C30C30C30C30C30C30C303C30C3C02A8" ;
	    attribute INITP_01 of bram : label is "EF0FAA2CCCCCCCCCCCECCCCCCCCCCCECCCECECCAC0A02C3E2A8B081330CC3333" ;
	    attribute INITP_02 of bram : label is "333333333332CCCCCCCCCCCCCCCBCCCCCCCCEDF333333B333333333CCCCCCCCC" ;
	    attribute INITP_03 of bram : label is "00000000000000000000000000000000000000C302FDD3267499D235C030CB33" ;
	    attribute INITP_04 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_05 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_06 of bram : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
	    attribute INITP_07 of bram : label is "C000000000000000000000000000000000000000000000000000000000000000" ;
	begin
	    bram : component RAMB16_S9_S18
	        generic map (
	            INIT_00 => X"BFE00F02147DBFE00F01C0010137020003000D000E00CF04CF01CF00CF070F00",
	            INIT_01 => X"1F705066EF481F70505FEF4C1F70505FEF6C1F70AEFD400B149ABFE00F041415",
	            INIT_02 => X"EF721F70504CEF531F70504CEF731F705047EF411F705047EF611F705066EF68",
	            INIT_03 => X"506BEF541F70506BEF741F70505BEF441F70505BEF641F705051EF521F705051",
	            INIT_04 => X"00B700BB13F00186A00000B700BB12F00186A000506FEF581F70506FEF781F70",
	            INIT_05 => X"0186A00000B700FF00BBA00000B700DB00A700A3CF040F01C202C30300BBA000",
	            INIT_06 => X"00BBA00000B7012600BBA00000B700BB11F00186A00000B700C300BBCE0410F0",
	            INIT_07 => X"DFF01FD0AEFEA000547ACF010F05A00000B70169CF070F000079CF070F01014A",
	            INIT_08 => X"1AC05491EF031FD0409219C0548CEF021FD0409218C05487EF01409217C05483",
	            INIT_09 => X"0F03C101C000C202C303AEFBA00000B70D00CE02B400FFC00F0D8D010DFF4092",
	            INIT_0A => X"54ADAF024F0414F0A000CF040F0041024001A00050A3AF014F0040A900A3CF04",
	            INIT_0B => X"00AC0F6B00AC0F4F00B2A00000AC0F3E00B2A00000AC0F0A00AC0F0DA000C405",
	            INIT_0C => X"00AC0F2000F31F0000F31F1000AC0F2000AC0F7200AC0F5700B2A00000AC0F21",
	            INIT_0D => X"00AC0F6400AC0F5200B2A00000F31F2000F31F3000AC0F2000AC0F7400AC0F61",
	            INIT_0E => X"00F31F3000AC0F2000AC0F7400AC0F6100AC0F2000F31F0000F31F1000AC0F20",
	            INIT_0F => X"00B2A00000AC019CAF0F1F5000AC019C0F0E0F0E0F0E0F0E15F0A00000F31F20",
	            INIT_10 => X"00F31F3000AC0F2000AC0F3D00AC0F2000AC0F7200AC0F6400AC0F6400AC0F41",
	            INIT_11 => X"0F2000AC0F3D00AC0F2000AC0F6100AC0F7400AC0F6100AC0F4400B200F31F20",
	            INIT_12 => X"0F7300AC0F6900AC0F2000AC1F9000AC1F8000B2A00000F31F0000F31F1000AC",
	            INIT_13 => X"00AC0F5200AC0F4500AC0F5000AC0F4100B2A00000AC8F30018600AC0F2000AC",
	            INIT_14 => X"00AC0F6600AC0F6F00AC0F53A00000B700AC0F3100AC0F3100AC0F2000AC0F54",
	            INIT_15 => X"00AC0F2000AC0F7400AC0F6500AC0F7300AC0F6500AC0F5200AC0F2000AC0F74",
	            INIT_16 => X"0F7400AC0F6600AC0F6F00AC0F53A00000AC0F6800AC0F6700AC0F6900AC0F48",
	            INIT_17 => X"0F4C00AC0F2000AC0F7400AC0F6500AC0F7300AC0F6500AC0F5200AC0F2000AC",
	            INIT_18 => X"5193B880A80FA90F19F001951F9018F001951F80A00000AC0F7700AC0F6F00AC",
	            INIT_19 => X"8F305DA1C40A14F0A000CF37A000CF305D9AC44014F0A0001F90418EC8018910",
	            INIT_1A => X"1FC04C0316F0A00000B700BB55A4850100AC8F301F5000B205EAA0008F37A000",
	            INIT_1B => X"00000000000000000000000000000000000000000000000080011F600E0100AC",
	            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INIT_3F => X"41AD000000000000000000000000000000000000000000000000000000000000",
	            INITP_00 => X"02D2F8E3EFEF3BF0EFEFF8AEF3BCEC30C30C30C30C30C30C30C303C30C3C02A8",
	            INITP_01 => X"EF0FAA2CCCCCCCCCCCECCCCCCCCCCCECCCECECCAC0A02C3E2A8B081330CC3333",
	            INITP_02 => X"333333333332CCCCCCCCCCCCCCCBCCCCCCCCEDF333333B333333333CCCCCCCCC",
	            INITP_03 => X"00000000000000000000000000000000000000C302FDD3267499D235C030CB33",
	            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
	            INITP_07 => X"C000000000000000000000000000000000000000000000000000000000000000"
	        )
	        port map (
	            DIB => "0000000000000000",
	            DIPB => "00",
	            ENB => '1',
	            WEB => '0',
	            SSRB => '0',
	            CLKB => clk,
	            ADDRB => address,
	            DOB => instruction( INSTSIZE - 3 downto 0 ),
	            DOPB => instruction( INSTSIZE - 1 downto INSTSIZE - 2 ),
	            DIA => jdata( JDATASIZE - 2 downto 0 ),
	            DIPA => jdata( JDATASIZE - 1 downto JDATASIZE - 1 ),
	            ENA => juser1,
	            WEA => jwrite,
	            SSRA => '0',
	            CLKA => clk,
	            ADDRA => jaddr,
	            DOA => open,
	            DOPA => open 
	        ) ;
	end generate ;

	I16 : if PicoType = pbtI generate
		attribute INIT_00 of bram : label is "BFE00F02147DBFE00F01C0010137020003000D000E00CF04CF01CF00CF070F00" ;
		attribute INIT_01 of bram : label is "1F705066EF481F70505FEF4C1F70505FEF6C1F70AEFD400B149ABFE00F041415" ;
		attribute INIT_02 of bram : label is "EF721F70504CEF531F70504CEF731F705047EF411F705047EF611F705066EF68" ;
		attribute INIT_03 of bram : label is "506BEF541F70506BEF741F70505BEF441F70505BEF641F705051EF521F705051" ;
		attribute INIT_04 of bram : label is "00B700BB13F00186A00000B700BB12F00186A000506FEF581F70506FEF781F70" ;
		attribute INIT_05 of bram : label is "0186A00000B700FF00BBA00000B700DB00A700A3CF040F01C202C30300BBA000" ;
		attribute INIT_06 of bram : label is "00BBA00000B7012600BBA00000B700BB11F00186A00000B700C300BBCE0410F0" ;
		attribute INIT_07 of bram : label is "DFF01FD0AEFEA000547ACF010F05A00000B70169CF070F000079CF070F01014A" ;
		attribute INIT_08 of bram : label is "1AC05491EF031FD0409219C0548CEF021FD0409218C05487EF01409217C05483" ;
		attribute INIT_09 of bram : label is "0F03C101C000C202C303AEFBA00000B70D00CE02B400FFC00F0D8D010DFF4092" ;
		attribute INIT_0A of bram : label is "54ADAF024F0414F0A000CF040F0041024001A00050A3AF014F0040A900A3CF04" ;
		attribute INIT_0B of bram : label is "00AC0F6B00AC0F4F00B2A00000AC0F3E00B2A00000AC0F0A00AC0F0DA000C405" ;
		attribute INIT_0C of bram : label is "00AC0F2000F31F0000F31F1000AC0F2000AC0F7200AC0F5700B2A00000AC0F21" ;
		attribute INIT_0D of bram : label is "00AC0F6400AC0F5200B2A00000F31F2000F31F3000AC0F2000AC0F7400AC0F61" ;
		attribute INIT_0E of bram : label is "00F31F3000AC0F2000AC0F7400AC0F6100AC0F2000F31F0000F31F1000AC0F20" ;
		attribute INIT_0F of bram : label is "00B2A00000AC019CAF0F1F5000AC019C0F0E0F0E0F0E0F0E15F0A00000F31F20" ;
	begin
	    bram : component RAMB4_S8_S16
	        generic map (
	            INIT_00 => X"BFE00F02147DBFE00F01C0010137020003000D000E00CF04CF01CF00CF070F00",
	            INIT_01 => X"1F705066EF481F70505FEF4C1F70505FEF6C1F70AEFD400B149ABFE00F041415",
	            INIT_02 => X"EF721F70504CEF531F70504CEF731F705047EF411F705047EF611F705066EF68",
	            INIT_03 => X"506BEF541F70506BEF741F70505BEF441F70505BEF641F705051EF521F705051",
	            INIT_04 => X"00B700BB13F00186A00000B700BB12F00186A000506FEF581F70506FEF781F70",
	            INIT_05 => X"0186A00000B700FF00BBA00000B700DB00A700A3CF040F01C202C30300BBA000",
	            INIT_06 => X"00BBA00000B7012600BBA00000B700BB11F00186A00000B700C300BBCE0410F0",
	            INIT_07 => X"DFF01FD0AEFEA000547ACF010F05A00000B70169CF070F000079CF070F01014A",
	            INIT_08 => X"1AC05491EF031FD0409219C0548CEF021FD0409218C05487EF01409217C05483",
	            INIT_09 => X"0F03C101C000C202C303AEFBA00000B70D00CE02B400FFC00F0D8D010DFF4092",
	            INIT_0A => X"54ADAF024F0414F0A000CF040F0041024001A00050A3AF014F0040A900A3CF04",
	            INIT_0B => X"00AC0F6B00AC0F4F00B2A00000AC0F3E00B2A00000AC0F0A00AC0F0DA000C405",
	            INIT_0C => X"00AC0F2000F31F0000F31F1000AC0F2000AC0F7200AC0F5700B2A00000AC0F21",
	            INIT_0D => X"00AC0F6400AC0F5200B2A00000F31F2000F31F3000AC0F2000AC0F7400AC0F61",
	            INIT_0E => X"00F31F3000AC0F2000AC0F7400AC0F6100AC0F2000F31F0000F31F1000AC0F20",
	            INIT_0F => X"00B2A00000AC019CAF0F1F5000AC019C0F0E0F0E0F0E0F0E15F0A00000F31F20"
	        )
			port map (
				DIB => "0000000000000000",  
				ENB => '1', 
				WEB => '0',
				RSTB =>	'0',
				CLKB => clk,
				ADDRB => address,
				DOB => instruction( INSTSIZE - 1 downto 0 ),  
				DIA => jdata( JDATASIZE - 1 downto 0 ),   
				ENA => juser1, 
				WEA => jwrite,
				RSTA => '0',
				CLKA => clk,
				ADDRA => jaddr,
				DOA => open  
			) ; 
	end generate ;

	I20 : if PicoType = pbtS generate
		attribute INIT_00 of ram_1 : label is "3003003003003003003003003003003003003003000330030030033000022220" ;
		attribute INIT_01 of ram_1 : label is "0002310233203203323332330323330032333233332022323303233032300300" ;
		attribute INIT_02 of ram_1 : label is "3030323032303022300022000230033202222023002001030300303003030303" ;
		attribute INIT_03 of ram_1 : label is "3233003322220230303030303030303030303230303030303030303030303230" ;
		attribute INIT_04 of ram_1 : label is "3030303032313303030303030323030303030303030303303030303030303030" ;
		attribute INIT_05 of ram_1 : label is "0303030303030303030303023030303030303030303030303030302330303030" ;
		attribute INIT_06 of ram_1 : label is "0000000000003003000233313103021213102121310203113000030030230303" ;
		attribute INIT_07 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_1 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_1 : label is "3000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_2 : label is "5E15E15E15E15E15E15E15E15E15E15E15E15E15E1A41B01B01B0C00000CCCC0" ;
		attribute INIT_01 of ram_2 : label is "D1AA5C0A00C00C000A000A0010A000C10A000A0000C0CC0A0010A0010A5E15E1" ;
		attribute INIT_02 of ram_2 : label is "00000A000A0000AC5A41AC044A5A440C0CCCCAA00CBF080415E1415E1415E415" ;
		attribute INIT_03 of ram_2 : label is "0A00A10000001A01010000000001010000000A01010000000001010000000A00" ;
		attribute INIT_04 of ram_2 : label is "000000000A0800000000001010A0101000000000000000010100000000000000" ;
		attribute INIT_05 of ram_2 : label is "00000000000000000000000A000000000000000000000000000000A000000000" ;
		attribute INIT_06 of ram_2 : label is "0000000000008100141A005808100A8A85C1ACAC5C1A14C85BAA101101A00000" ;
		attribute INIT_07 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_2 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_2 : label is "4000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_3 : label is "0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FFE04FF4FF4FF0123DEFFFFF" ;
		attribute INIT_01 of ram_3 : label is "FFE04FF001FF0FF100010000110000E01000000000FF230000310002100FF0FF" ;
		attribute INIT_02 of ram_3 : label is "0F0F000F000F0F044FF40FF1000FF00FF1023E00DE4FFDD0A4FF094FF084F074" ;
		attribute INIT_03 of ram_3 : label is "0001FF01FFFF500F0F0F0F0F0F0F0F0F0F0F000F0F0F0F0F0F0F0F0F0F0F000F" ;
		attribute INIT_04 of ram_3 : label is "0F0F0F0F000F10F0F0F0F0F0F000F0F0F0F0F0F0F0F0F00F0F0F0F0F0F0F0F0F" ;
		attribute INIT_05 of ram_3 : label is "F0F0F0F0F0F0F0F0F0F0F0F00F0F0F0F0F0F0F0F0F0F0F0F0F0F0F000F0F0F0F" ;
		attribute INIT_06 of ram_3 : label is "0000000000000FE0FC6000550FF050F0FD440F0FD440F189188991F81F00F0F0" ;
		attribute INIT_07 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_3 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_3 : label is "1000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_4 : label is "657677547567557577457477447467667647547567F09E01E07E003000000000" ;
		attribute INIT_01 of ram_4 : label is "FDF07000B6007004B0B2B0BBF80BCB0F80BFB0BDAA0000B0BBF80BBF80657677" ;
		attribute INIT_02 of ram_4 : label is "A6A4B0A3B0A0A000A00F000000A00AA000000F0B000C00F9C90D9C80D9C809C8" ;
		attribute INIT_03 of ram_4 : label is "B0A905A90000F0F2F3A2A7A6A2F0F1A2A6A5B0F2F3A2A7A6A2F0F1A2A7A5B0A2" ;
		attribute INIT_04 of ram_4 : label is "A5A4A5A4B0A38A2A7A6A2A9A8B0F0F1A2A3A2A6A7A6A4BF2F3A2A3A2A7A6A6A4" ;
		attribute INIT_05 of ram_4 : label is "4A2A7A6A7A6A5A2A7A6A6A50A6A6A6A4A2A7A6A7A6A5A2A7A6A6A50BA3A3A2A5" ;
		attribute INIT_06 of ram_4 : label is "000000000000060AC0F0BBA0A35BE0303A0F030394F098019800F99F980A7A6A" ;
		attribute INIT_07 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_4 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_4 : label is "A000000000000000000000000000000000000000000000000000000000000000" ;

		attribute INIT_00 of ram_5 : label is "B40B40B40B40120120C30C30710710680680FC0FC0DBA04502D0117000041070" ;
		attribute INIT_01 of ram_5 : label is "00E0A1507970971AB076B07B06073B40607FB07B734123B07B0607B060F80F80" ;
		attribute INIT_02 of ram_5 : label is "CBCF20CE20CACD05D24004021031093431023B070200D1F2013020C202071203" ;
		attribute INIT_03 of ram_5 : label is "20CCF0CCEEEE003030C0C4C1C03030C0C4C2203030C0C4C1C03030C0C2C720C1" ;
		attribute INIT_04 of ram_5 : label is "C2C5C0C120C06C0C3C9C0C0C0203030C0CDC0C1C4C1C423030C0CDC0C2C4C4C1" ;
		attribute INIT_05 of ram_5 : label is "CC0C4C5C3C5C2C0C4C6CFC30C8C7C9C8C0C4C5C3C5C2C0C4C6CFC307C1C1C0C4" ;
		attribute INIT_06 of ram_5 : label is "000000000000101C03007B41C002A07001A00700A0000E1030FF0500500C7CFC" ;
		attribute INIT_07 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_08 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_09 of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0A of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0B of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0C of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0D of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0E of ram_5 : label is "0000000000000000000000000000000000000000000000000000000000000000" ;
		attribute INIT_0F of ram_5 : label is "D000000000000000000000000000000000000000000000000000000000000000" ;

		signal data_out : std_logic_vector( 3 downto 0 ) ;
	begin
	    ram_1 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"3003003003003003003003003003003003003003000330030030033000022220",
				INIT_01 => X"0002310233203203323332330323330032333233332022323303233032300300",
				INIT_02 => X"3030323032303022300022000230033202222023002001030300303003030303",
				INIT_03 => X"3233003322220230303030303030303030303230303030303030303030303230",
				INIT_04 => X"3030303032313303030303030323030303030303030303303030303030303030",
				INIT_05 => X"0303030303030303030303023030303030303030303030303030302330303030",
				INIT_06 => X"0000000000003003000233313103021213102121310203113000030030230303",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"3000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => data_out,  
				DIB => jdata( JDATASIZE - 1 downto 16 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
			-- loose top 2 bits
			instruction( 17 downto 16 ) <= data_out( 1 downto 0 ) ;

	    ram_2 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"5E15E15E15E15E15E15E15E15E15E15E15E15E15E1A41B01B01B0C00000CCCC0",
				INIT_01 => X"D1AA5C0A00C00C000A000A0010A000C10A000A0000C0CC0A0010A0010A5E15E1",
				INIT_02 => X"00000A000A0000AC5A41AC044A5A440C0CCCCAA00CBF080415E1415E1415E415",
				INIT_03 => X"0A00A10000001A01010000000001010000000A01010000000001010000000A00",
				INIT_04 => X"000000000A0800000000001010A0101000000000000000010100000000000000",
				INIT_05 => X"00000000000000000000000A000000000000000000000000000000A000000000",
				INIT_06 => X"0000000000008100141A005808100A8A85C1ACAC5C1A14C85BAA101101A00000",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"4000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 15 downto 12 ),  
				DIB => jdata( 15 downto 12 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_3 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FF0FFE04FF4FF4FF0123DEFFFFF",
				INIT_01 => X"FFE04FF001FF0FF100010000110000E01000000000FF230000310002100FF0FF",
				INIT_02 => X"0F0F000F000F0F044FF40FF1000FF00FF1023E00DE4FFDD0A4FF094FF084F074",
				INIT_03 => X"0001FF01FFFF500F0F0F0F0F0F0F0F0F0F0F000F0F0F0F0F0F0F0F0F0F0F000F",
				INIT_04 => X"0F0F0F0F000F10F0F0F0F0F0F000F0F0F0F0F0F0F0F0F00F0F0F0F0F0F0F0F0F",
				INIT_05 => X"F0F0F0F0F0F0F0F0F0F0F0F00F0F0F0F0F0F0F0F0F0F0F0F0F0F0F000F0F0F0F",
				INIT_06 => X"0000000000000FE0FC6000550FF050F0FD440F0FD440F189188991F81F00F0F0",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"1000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 11 downto 8 ),  
				DIB => jdata( 11 downto 8 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_4 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"657677547567557577457477447467667647547567F09E01E07E003000000000",
				INIT_01 => X"FDF07000B6007004B0B2B0BBF80BCB0F80BFB0BDAA0000B0BBF80BBF80657677",
				INIT_02 => X"A6A4B0A3B0A0A000A00F000000A00AA000000F0B000C00F9C90D9C80D9C809C8",
				INIT_03 => X"B0A905A90000F0F2F3A2A7A6A2F0F1A2A6A5B0F2F3A2A7A6A2F0F1A2A7A5B0A2",
				INIT_04 => X"A5A4A5A4B0A38A2A7A6A2A9A8B0F0F1A2A3A2A6A7A6A4BF2F3A2A3A2A7A6A6A4",
				INIT_05 => X"4A2A7A6A7A6A5A2A7A6A6A50A6A6A6A4A2A7A6A7A6A5A2A7A6A6A50BA3A3A2A5",
				INIT_06 => X"000000000000060AC0F0BBA0A35BE0303A0F030394F098019800F99F980A7A6A",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"A000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 7 downto 4 ),  
				DIB => jdata( 7 downto 4 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 

	    ram_5 : component RAMB4_S4_S4
	        generic map (
				INIT_00 => X"B40B40B40B40120120C30C30710710680680FC0FC0DBA04502D0117000041070",
				INIT_01 => X"00E0A1507970971AB076B07B06073B40607FB07B734123B07B0607B060F80F80",
				INIT_02 => X"CBCF20CE20CACD05D24004021031093431023B070200D1F2013020C202071203",
				INIT_03 => X"20CCF0CCEEEE003030C0C4C1C03030C0C4C2203030C0C4C1C03030C0C2C720C1",
				INIT_04 => X"C2C5C0C120C06C0C3C9C0C0C0203030C0CDC0C1C4C1C423030C0CDC0C2C4C4C1",
				INIT_05 => X"CC0C4C5C3C5C2C0C4C6CFC30C8C7C9C8C0C4C5C3C5C2C0C4C6CFC307C1C1C0C4",
				INIT_06 => X"000000000000101C03007B41C002A07001A00700A0000E1030FF0500500C7CFC",
				INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
				INIT_0F => X"D000000000000000000000000000000000000000000000000000000000000000"
	        )
			port map (
				DIA => "0000",  
				ENA => '1', 
				WEA => '0',
				RSTA =>	'0',
				CLKA => clk,
				ADDRA => address,
				DOA => instruction( 3 downto 0 ),  
				DIB => jdata( 3 downto 0 ),   
				ENB => juser1, 
				WEB => jwrite,
				RSTB => '0',
				CLKB => clk,
				ADDRB => jaddr,
				DOB => open  
			) ; 
	end generate ;

	jdata <= ( others => '0' ) ;
	jaddr <= ( others => '0' ) ;
	juser1 <= '0' ;
	jwrite <= '0' ;
end architecture mix ;
